`timescale 1 ns / 10ps

//////////////////////////////////////////////////////////////////////////////////
// Company: Fudan University
// Engineer: CaiChang
// 
// Create Date: 2021/12/01 11:00:11
// Design Name: 
// Module Name: wallace_tree
// Project Name: multiplier
// Target Devices: 
// Tool Versions: 
// Description: 
//              a 32x32 multiplier with booth2 algorithm and jump wallace tree
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////\

module wallace_tree(
    input [32 : 0] p0,
    input [32 : 0] p1,
    input [32 : 0] p2,
    input [32 : 0] p3,
    input [32 : 0] p4,
    input [32 : 0] p5,
    input [32 : 0] p6,
    input [32 : 0] p7,
    input [32 : 0] p8,
    input [32 : 0] p9,
    input [32 : 0] p10,
    input [32 : 0] p11,
    input [32 : 0] p12,
    input [32 : 0] p13,
    input [32 : 0] p14,
    input [32 : 0] p15,
    input [15 : 0] E,
    input [31 : 0] y,
    output [63 : 0] add0,
    output [63 : 0] add1
);

wire [34 : 0] CSA0_s,CSA0_co;
wire [34 : 0] CSA1_s,CSA1_co;
wire [34 : 0] CSA2_s,CSA2_co;
wire [34 : 0] CSA3_s,CSA3_co;
wire [34 : 0] CSA4_s,CSA4_co;
wire [33 : 0] com_s;
wire [33 : 0] com_co;
wire [25 : 0] com_ca;
wire [16 : 0] CSA5_s,CSA5_co;
wire [32 : 0] CSA6_s,CSA6_co;
wire [34 : 0] CSA7_s,CSA7_co;
wire [49 : 0] CSA8_s,CSA8_co;
wire [27 : 0] CSA9_s,CSA9_co;
wire [46 : 0] CSA10_s,CSA10_co;
wire [44 : 0] CSA11_s,CSA11_co;




//CSA0
fa CSA0_0
(
    .a(p0[2]),
    .b(p1[0]),
    .c(y[3]),
    .s(CSA0_s[0]),
    .co(CSA0_co[0])
);
ha CSA0_1
(
    .a(p0[3]),
    .b(p1[1]),
    .s(CSA0_s[1]),
    .co(CSA0_co[1])
);
fa CSA0_2
(
    .a(p0[4]),
    .b(p1[2]),
    .c(p2[0]),
    .s(CSA0_s[2]),
    .co(CSA0_co[2])
);
fa CSA0_3
(
    .a(p0[5]),
    .b(p1[3]),
    .c(p2[1]),
    .s(CSA0_s[3]),
    .co(CSA0_co[3])
);
fa CSA0_4
(
    .a(p0[6]),
    .b(p1[4]),
    .c(p2[2]),
    .s(CSA0_s[4]),
    .co(CSA0_co[4])
);
fa CSA0_5
(
    .a(p0[7]),
    .b(p1[5]),
    .c(p2[3]),
    .s(CSA0_s[5]),
    .co(CSA0_co[5])
);
fa CSA0_6
(
    .a(p0[8]),
    .b(p1[6]),
    .c(p2[4]),
    .s(CSA0_s[6]),
    .co(CSA0_co[6])
);
fa CSA0_7
(
    .a(p0[9]),
    .b(p1[7]),
    .c(p2[5]),
    .s(CSA0_s[7]),
    .co(CSA0_co[7])
);
fa CSA0_8
(
    .a(p0[10]),
    .b(p1[8]),
    .c(p2[6]),
    .s(CSA0_s[8]),
    .co(CSA0_co[8])
);
fa CSA0_9
(
    .a(p0[11]),
    .b(p1[9]),
    .c(p2[7]),
    .s(CSA0_s[9]),
    .co(CSA0_co[9])
);
fa CSA0_10
(
    .a(p0[12]),
    .b(p1[10]),
    .c(p2[8]),
    .s(CSA0_s[10]),
    .co(CSA0_co[10])
);
fa CSA0_11
(
    .a(p0[13]),
    .b(p1[11]),
    .c(p2[9]),
    .s(CSA0_s[11]),
    .co(CSA0_co[11])
);
fa CSA0_12
(
    .a(p0[14]),
    .b(p1[12]),
    .c(p2[10]),
    .s(CSA0_s[12]),
    .co(CSA0_co[12])
);
fa CSA0_13
(
    .a(p0[15]),
    .b(p1[13]),
    .c(p2[11]),
    .s(CSA0_s[13]),
    .co(CSA0_co[13])
);
fa CSA0_14
(
    .a(p0[16]),
    .b(p1[14]),
    .c(p2[12]),
    .s(CSA0_s[14]),
    .co(CSA0_co[14])
);
fa CSA0_15
(
    .a(p0[17]),
    .b(p1[15]),
    .c(p2[13]),
    .s(CSA0_s[15]),
    .co(CSA0_co[15])
);
fa CSA0_16
(
    .a(p0[18]),
    .b(p1[16]),
    .c(p2[14]),
    .s(CSA0_s[16]),
    .co(CSA0_co[16])
);
fa CSA0_17
(
    .a(p0[19]),
    .b(p1[17]),
    .c(p2[15]),
    .s(CSA0_s[17]),
    .co(CSA0_co[17])
);
fa CSA0_18
(
    .a(p0[20]),
    .b(p1[18]),
    .c(p2[16]),
    .s(CSA0_s[18]),
    .co(CSA0_co[18])
);
fa CSA0_19
(
    .a(p0[21]),
    .b(p1[19]),
    .c(p2[17]),
    .s(CSA0_s[19]),
    .co(CSA0_co[19])
);
fa CSA0_20
(
    .a(p0[22]),
    .b(p1[20]),
    .c(p2[18]),
    .s(CSA0_s[20]),
    .co(CSA0_co[20])
);
fa CSA0_21
(
    .a(p0[23]),
    .b(p1[21]),
    .c(p2[19]),
    .s(CSA0_s[21]),
    .co(CSA0_co[21])
);
fa CSA0_22
(
    .a(p0[24]),
    .b(p1[22]),
    .c(p2[20]),
    .s(CSA0_s[22]),
    .co(CSA0_co[22])
);
fa CSA0_23
(
    .a(p0[25]),
    .b(p1[23]),
    .c(p2[21]),
    .s(CSA0_s[23]),
    .co(CSA0_co[23])
);
fa CSA0_24
(
    .a(p0[26]),
    .b(p1[24]),
    .c(p2[22]),
    .s(CSA0_s[24]),
    .co(CSA0_co[24])
);
fa CSA0_25
(
    .a(p0[27]),
    .b(p1[25]),
    .c(p2[23]),
    .s(CSA0_s[25]),
    .co(CSA0_co[25])
);
fa CSA0_26
(
    .a(p0[28]),
    .b(p1[26]),
    .c(p2[24]),
    .s(CSA0_s[26]),
    .co(CSA0_co[26])
);
fa CSA0_27
(
    .a(p0[29]),
    .b(p1[27]),
    .c(p2[25]),
    .s(CSA0_s[27]),
    .co(CSA0_co[27])
);
fa CSA0_28
(
    .a(p0[30]),
    .b(p1[28]),
    .c(p2[26]),
    .s(CSA0_s[28]),
    .co(CSA0_co[28])
);
fa CSA0_29
(
    .a(p0[31]),
    .b(p1[29]),
    .c(p2[27]),
    .s(CSA0_s[29]),
    .co(CSA0_co[29])
);
fa CSA0_30
(
    .a(p0[32]),
    .b(p1[30]),
    .c(p2[28]),
    .s(CSA0_s[30]),
    .co(CSA0_co[30])
);
fa CSA0_31
(
    .a(~E[0]),
    .b(p1[31]),
    .c(p2[29]),
    .s(CSA0_s[31]),
    .co(CSA0_co[31])
);
fa CSA0_32
(
    .a(~E[0]),
    .b(p1[32]),
    .c(p2[30]),
    .s(CSA0_s[32]),
    .co(CSA0_co[32])
);
fa CSA0_33
(
    .a(E[0]),
    .b(E[1]),
    .c(p2[31]),
    .s(CSA0_s[33]),
    .co(CSA0_co[33])
);
ha CSA0_34
(
    .a(1'b1),
    .b(p2[32]),
    .s(CSA0_s[34]),
    .co(CSA0_co[34])
);

//CSA1
fa CSA1_0
(
    .a(p3[2]),
    .b(p4[0]),
    .c(y[9]),
    .s(CSA1_s[0]),
    .co(CSA1_co[0])
);
ha CSA1_1
(
    .a(p3[3]),
    .b(p4[1]),
    .s(CSA1_s[1]),
    .co(CSA1_co[1])
);
fa CSA1_2
(
    .a(p3[4]),
    .b(p4[2]),
    .c(p5[0]),
    .s(CSA1_s[2]),
    .co(CSA1_co[2])
);
fa CSA1_3
(
    .a(p3[5]),
    .b(p4[3]),
    .c(p5[1]),
    .s(CSA1_s[3]),
    .co(CSA1_co[3])
);
fa CSA1_4
(
    .a(p3[6]),
    .b(p4[4]),
    .c(p5[2]),
    .s(CSA1_s[4]),
    .co(CSA1_co[4])
);
fa CSA1_5
(
    .a(p3[7]),
    .b(p4[5]),
    .c(p5[3]),
    .s(CSA1_s[5]),
    .co(CSA1_co[5])
);
fa CSA1_6
(
    .a(p3[8]),
    .b(p4[6]),
    .c(p5[4]),
    .s(CSA1_s[6]),
    .co(CSA1_co[6])
);
fa CSA1_7
(
    .a(p3[9]),
    .b(p4[7]),
    .c(p5[5]),
    .s(CSA1_s[7]),
    .co(CSA1_co[7])
);
fa CSA1_8
(
    .a(p3[10]),
    .b(p4[8]),
    .c(p5[6]),
    .s(CSA1_s[8]),
    .co(CSA1_co[8])
);
fa CSA1_9
(
    .a(p3[11]),
    .b(p4[9]),
    .c(p5[7]),
    .s(CSA1_s[9]),
    .co(CSA1_co[9])
);
fa CSA1_10
(
    .a(p3[12]),
    .b(p4[10]),
    .c(p5[8]),
    .s(CSA1_s[10]),
    .co(CSA1_co[10])
);
fa CSA1_11
(
    .a(p3[13]),
    .b(p4[11]),
    .c(p5[9]),
    .s(CSA1_s[11]),
    .co(CSA1_co[11])
);
fa CSA1_12
(
    .a(p3[14]),
    .b(p4[12]),
    .c(p5[10]),
    .s(CSA1_s[12]),
    .co(CSA1_co[12])
);
fa CSA1_13
(
    .a(p3[15]),
    .b(p4[13]),
    .c(p5[11]),
    .s(CSA1_s[13]),
    .co(CSA1_co[13])
);
fa CSA1_14
(
    .a(p3[16]),
    .b(p4[14]),
    .c(p5[12]),
    .s(CSA1_s[14]),
    .co(CSA1_co[14])
);
fa CSA1_15
(
    .a(p3[17]),
    .b(p4[15]),
    .c(p5[13]),
    .s(CSA1_s[15]),
    .co(CSA1_co[15])
);
fa CSA1_16
(
    .a(p3[18]),
    .b(p4[16]),
    .c(p5[14]),
    .s(CSA1_s[16]),
    .co(CSA1_co[16])
);
fa CSA1_17
(
    .a(p3[19]),
    .b(p4[17]),
    .c(p5[15]),
    .s(CSA1_s[17]),
    .co(CSA1_co[17])
);
fa CSA1_18
(
    .a(p3[20]),
    .b(p4[18]),
    .c(p5[16]),
    .s(CSA1_s[18]),
    .co(CSA1_co[18])
);
fa CSA1_19
(
    .a(p3[21]),
    .b(p4[19]),
    .c(p5[17]),
    .s(CSA1_s[19]),
    .co(CSA1_co[19])
);
fa CSA1_20
(
    .a(p3[22]),
    .b(p4[20]),
    .c(p5[18]),
    .s(CSA1_s[20]),
    .co(CSA1_co[20])
);
fa CSA1_21
(
    .a(p3[23]),
    .b(p4[21]),
    .c(p5[19]),
    .s(CSA1_s[21]),
    .co(CSA1_co[21])
);
fa CSA1_22
(
    .a(p3[24]),
    .b(p4[22]),
    .c(p5[20]),
    .s(CSA1_s[22]),
    .co(CSA1_co[22])
);
fa CSA1_23
(
    .a(p3[25]),
    .b(p4[23]),
    .c(p5[21]),
    .s(CSA1_s[23]),
    .co(CSA1_co[23])
);
fa CSA1_24
(
    .a(p3[26]),
    .b(p4[24]),
    .c(p5[22]),
    .s(CSA1_s[24]),
    .co(CSA1_co[24])
);
fa CSA1_25
(
    .a(p3[27]),
    .b(p4[25]),
    .c(p5[23]),
    .s(CSA1_s[25]),
    .co(CSA1_co[25])
);
fa CSA1_26
(
    .a(p3[28]),
    .b(p4[26]),
    .c(p5[24]),
    .s(CSA1_s[26]),
    .co(CSA1_co[26])
);
fa CSA1_27
(
    .a(p3[29]),
    .b(p4[27]),
    .c(p5[25]),
    .s(CSA1_s[27]),
    .co(CSA1_co[27])
);
fa CSA1_28
(
    .a(p3[30]),
    .b(p4[28]),
    .c(p5[26]),
    .s(CSA1_s[28]),
    .co(CSA1_co[28])
);
fa CSA1_29
(
    .a(p3[31]),
    .b(p4[29]),
    .c(p5[27]),
    .s(CSA1_s[29]),
    .co(CSA1_co[29])
);
fa CSA1_30
(
    .a(p3[32]),
    .b(p4[30]),
    .c(p5[28]),
    .s(CSA1_s[30]),
    .co(CSA1_co[30])
);
fa CSA1_31
(
    .a(E[3]),
    .b(p4[31]),
    .c(p5[29]),
    .s(CSA1_s[31]),
    .co(CSA1_co[31])
);
fa CSA1_32
(
    .a(1'b1),
    .b(p4[32]),
    .c(p5[30]),
    .s(CSA1_s[32]),
    .co(CSA1_co[32])
);
ha CSA1_33
(
    .a(E[4]),
    .b(p5[31]),
    .s(CSA1_s[33]),
    .co(CSA1_co[33])
);
ha CSA1_34
(
    .a(1'b1),
    .b(p5[32]),
    .s(CSA1_s[34]),
    .co(CSA1_co[34])
);

//CSA2
fa CSA2_0
(
    .a(p6[2]),
    .b(p7[0]),
    .c(y[15]),
    .s(CSA2_s[0]),
    .co(CSA2_co[0])
);
ha CSA2_1
(
    .a(p6[3]),
    .b(p7[1]),
    .s(CSA2_s[1]),
    .co(CSA2_co[1])
);
fa CSA2_2
(
    .a(p6[4]),
    .b(p7[2]),
    .c(p8[0]),
    .s(CSA2_s[2]),
    .co(CSA2_co[2])
);
fa CSA2_3
(
    .a(p6[5]),
    .b(p7[3]),
    .c(p8[1]),
    .s(CSA2_s[3]),
    .co(CSA2_co[3])
);
fa CSA2_4
(
    .a(p6[6]),
    .b(p7[4]),
    .c(p8[2]),
    .s(CSA2_s[4]),
    .co(CSA2_co[4])
);
fa CSA2_5
(
    .a(p6[7]),
    .b(p7[5]),
    .c(p8[3]),
    .s(CSA2_s[5]),
    .co(CSA2_co[5])
);
fa CSA2_6
(
    .a(p6[8]),
    .b(p7[6]),
    .c(p8[4]),
    .s(CSA2_s[6]),
    .co(CSA2_co[6])
);
fa CSA2_7
(
    .a(p6[9]),
    .b(p7[7]),
    .c(p8[5]),
    .s(CSA2_s[7]),
    .co(CSA2_co[7])
);
fa CSA2_8
(
    .a(p6[10]),
    .b(p7[8]),
    .c(p8[6]),
    .s(CSA2_s[8]),
    .co(CSA2_co[8])
);
fa CSA2_9
(
    .a(p6[11]),
    .b(p7[9]),
    .c(p8[7]),
    .s(CSA2_s[9]),
    .co(CSA2_co[9])
);
fa CSA2_10
(
    .a(p6[12]),
    .b(p7[10]),
    .c(p8[8]),
    .s(CSA2_s[10]),
    .co(CSA2_co[10])
);
fa CSA2_11
(
    .a(p6[13]),
    .b(p7[11]),
    .c(p8[9]),
    .s(CSA2_s[11]),
    .co(CSA2_co[11])
);
fa CSA2_12
(
    .a(p6[14]),
    .b(p7[12]),
    .c(p8[10]),
    .s(CSA2_s[12]),
    .co(CSA2_co[12])
);
fa CSA2_13
(
    .a(p6[15]),
    .b(p7[13]),
    .c(p8[11]),
    .s(CSA2_s[13]),
    .co(CSA2_co[13])
);
fa CSA2_14
(
    .a(p6[16]),
    .b(p7[14]),
    .c(p8[12]),
    .s(CSA2_s[14]),
    .co(CSA2_co[14])
);
fa CSA2_15
(
    .a(p6[17]),
    .b(p7[15]),
    .c(p8[13]),
    .s(CSA2_s[15]),
    .co(CSA2_co[15])
);
fa CSA2_16
(
    .a(p6[18]),
    .b(p7[16]),
    .c(p8[14]),
    .s(CSA2_s[16]),
    .co(CSA2_co[16])
);
fa CSA2_17
(
    .a(p6[19]),
    .b(p7[17]),
    .c(p8[15]),
    .s(CSA2_s[17]),
    .co(CSA2_co[17])
);
fa CSA2_18
(
    .a(p6[20]),
    .b(p7[18]),
    .c(p8[16]),
    .s(CSA2_s[18]),
    .co(CSA2_co[18])
);
fa CSA2_19
(
    .a(p6[21]),
    .b(p7[19]),
    .c(p8[17]),
    .s(CSA2_s[19]),
    .co(CSA2_co[19])
);
fa CSA2_20
(
    .a(p6[22]),
    .b(p7[20]),
    .c(p8[18]),
    .s(CSA2_s[20]),
    .co(CSA2_co[20])
);
fa CSA2_21
(
    .a(p6[23]),
    .b(p7[21]),
    .c(p8[19]),
    .s(CSA2_s[21]),
    .co(CSA2_co[21])
);
fa CSA2_22
(
    .a(p6[24]),
    .b(p7[22]),
    .c(p8[20]),
    .s(CSA2_s[22]),
    .co(CSA2_co[22])
);
fa CSA2_23
(
    .a(p6[25]),
    .b(p7[23]),
    .c(p8[21]),
    .s(CSA2_s[23]),
    .co(CSA2_co[23])
);
fa CSA2_24
(
    .a(p6[26]),
    .b(p7[24]),
    .c(p8[22]),
    .s(CSA2_s[24]),
    .co(CSA2_co[24])
);
fa CSA2_25
(
    .a(p6[27]),
    .b(p7[25]),
    .c(p8[23]),
    .s(CSA2_s[25]),
    .co(CSA2_co[25])
);
fa CSA2_26
(
    .a(p6[28]),
    .b(p7[26]),
    .c(p8[24]),
    .s(CSA2_s[26]),
    .co(CSA2_co[26])
);
fa CSA2_27
(
    .a(p6[29]),
    .b(p7[27]),
    .c(p8[25]),
    .s(CSA2_s[27]),
    .co(CSA2_co[27])
);
fa CSA2_28
(
    .a(p6[30]),
    .b(p7[28]),
    .c(p8[26]),
    .s(CSA2_s[28]),
    .co(CSA2_co[28])
);
fa CSA2_29
(
    .a(p6[31]),
    .b(p7[29]),
    .c(p8[27]),
    .s(CSA2_s[29]),
    .co(CSA2_co[29])
);
fa CSA2_30
(
    .a(p6[32]),
    .b(p7[30]),
    .c(p8[28]),
    .s(CSA2_s[30]),
    .co(CSA2_co[30])
);
fa CSA2_31
(
    .a(E[6]),
    .b(p7[31]),
    .c(p8[29]),
    .s(CSA2_s[31]),
    .co(CSA2_co[31])
);
fa CSA2_32
(
    .a(1'b1),
    .b(p7[32]),
    .c(p8[30]),
    .s(CSA2_s[32]),
    .co(CSA2_co[32])
);
ha CSA2_33
(
    .a(E[7]),
    .b(p8[31]),
    .s(CSA2_s[33]),
    .co(CSA2_co[33])
);
ha CSA2_34
(
    .a(1'b1),
    .b(p8[32]),
    .s(CSA2_s[34]),
    .co(CSA2_co[34])
);

//CSA3
fa CSA3_0
(
    .a(p9[2]),
    .b(p10[0]),
    .c(y[21]),
    .s(CSA3_s[0]),
    .co(CSA3_co[0])
);
ha CSA3_1
(
    .a(p9[3]),
    .b(p10[1]),
    .s(CSA3_s[1]),
    .co(CSA3_co[1])
);
fa CSA3_2
(
    .a(p9[4]),
    .b(p10[2]),
    .c(p11[0]),
    .s(CSA3_s[2]),
    .co(CSA3_co[2])
);
fa CSA3_3
(
    .a(p9[5]),
    .b(p10[3]),
    .c(p11[1]),
    .s(CSA3_s[3]),
    .co(CSA3_co[3])
);
fa CSA3_4
(
    .a(p9[6]),
    .b(p10[4]),
    .c(p11[2]),
    .s(CSA3_s[4]),
    .co(CSA3_co[4])
);
fa CSA3_5
(
    .a(p9[7]),
    .b(p10[5]),
    .c(p11[3]),
    .s(CSA3_s[5]),
    .co(CSA3_co[5])
);
fa CSA3_6
(
    .a(p9[8]),
    .b(p10[6]),
    .c(p11[4]),
    .s(CSA3_s[6]),
    .co(CSA3_co[6])
);
fa CSA3_7
(
    .a(p9[9]),
    .b(p10[7]),
    .c(p11[5]),
    .s(CSA3_s[7]),
    .co(CSA3_co[7])
);
fa CSA3_8
(
    .a(p9[10]),
    .b(p10[8]),
    .c(p11[6]),
    .s(CSA3_s[8]),
    .co(CSA3_co[8])
);
fa CSA3_9
(
    .a(p9[11]),
    .b(p10[9]),
    .c(p11[7]),
    .s(CSA3_s[9]),
    .co(CSA3_co[9])
);
fa CSA3_10
(
    .a(p9[12]),
    .b(p10[10]),
    .c(p11[8]),
    .s(CSA3_s[10]),
    .co(CSA3_co[10])
);
fa CSA3_11
(
    .a(p9[13]),
    .b(p10[11]),
    .c(p11[9]),
    .s(CSA3_s[11]),
    .co(CSA3_co[11])
);
fa CSA3_12
(
    .a(p9[14]),
    .b(p10[12]),
    .c(p11[10]),
    .s(CSA3_s[12]),
    .co(CSA3_co[12])
);
fa CSA3_13
(
    .a(p9[15]),
    .b(p10[13]),
    .c(p11[11]),
    .s(CSA3_s[13]),
    .co(CSA3_co[13])
);
fa CSA3_14
(
    .a(p9[16]),
    .b(p10[14]),
    .c(p11[12]),
    .s(CSA3_s[14]),
    .co(CSA3_co[14])
);
fa CSA3_15
(
    .a(p9[17]),
    .b(p10[15]),
    .c(p11[13]),
    .s(CSA3_s[15]),
    .co(CSA3_co[15])
);
fa CSA3_16
(
    .a(p9[18]),
    .b(p10[16]),
    .c(p11[14]),
    .s(CSA3_s[16]),
    .co(CSA3_co[16])
);
fa CSA3_17
(
    .a(p9[19]),
    .b(p10[17]),
    .c(p11[15]),
    .s(CSA3_s[17]),
    .co(CSA3_co[17])
);
fa CSA3_18
(
    .a(p9[20]),
    .b(p10[18]),
    .c(p11[16]),
    .s(CSA3_s[18]),
    .co(CSA3_co[18])
);
fa CSA3_19
(
    .a(p9[21]),
    .b(p10[19]),
    .c(p11[17]),
    .s(CSA3_s[19]),
    .co(CSA3_co[19])
);
fa CSA3_20
(
    .a(p9[22]),
    .b(p10[20]),
    .c(p11[18]),
    .s(CSA3_s[20]),
    .co(CSA3_co[20])
);
fa CSA3_21
(
    .a(p9[23]),
    .b(p10[21]),
    .c(p11[19]),
    .s(CSA3_s[21]),
    .co(CSA3_co[21])
);
fa CSA3_22
(
    .a(p9[24]),
    .b(p10[22]),
    .c(p11[20]),
    .s(CSA3_s[22]),
    .co(CSA3_co[22])
);
fa CSA3_23
(
    .a(p9[25]),
    .b(p10[23]),
    .c(p11[21]),
    .s(CSA3_s[23]),
    .co(CSA3_co[23])
);
fa CSA3_24
(
    .a(p9[26]),
    .b(p10[24]),
    .c(p11[22]),
    .s(CSA3_s[24]),
    .co(CSA3_co[24])
);
fa CSA3_25
(
    .a(p9[27]),
    .b(p10[25]),
    .c(p11[23]),
    .s(CSA3_s[25]),
    .co(CSA3_co[25])
);
fa CSA3_26
(
    .a(p9[28]),
    .b(p10[26]),
    .c(p11[24]),
    .s(CSA3_s[26]),
    .co(CSA3_co[26])
);
fa CSA3_27
(
    .a(p9[29]),
    .b(p10[27]),
    .c(p11[25]),
    .s(CSA3_s[27]),
    .co(CSA3_co[27])
);
fa CSA3_28
(
    .a(p9[30]),
    .b(p10[28]),
    .c(p11[26]),
    .s(CSA3_s[28]),
    .co(CSA3_co[28])
);
fa CSA3_29
(
    .a(p9[31]),
    .b(p10[29]),
    .c(p11[27]),
    .s(CSA3_s[29]),
    .co(CSA3_co[29])
);
fa CSA3_30
(
    .a(p9[32]),
    .b(p10[30]),
    .c(p11[28]),
    .s(CSA3_s[30]),
    .co(CSA3_co[30])
);
fa CSA3_31
(
    .a(E[9]),
    .b(p10[31]),
    .c(p11[29]),
    .s(CSA3_s[31]),
    .co(CSA3_co[31])
);
fa CSA3_32
(
    .a(1'b1),
    .b(p10[32]),
    .c(p11[30]),
    .s(CSA3_s[32]),
    .co(CSA3_co[32])
);
ha CSA3_33
(
    .a(E[10]),
    .b(p11[31]),
    .s(CSA3_s[33]),
    .co(CSA3_co[33])
);
ha CSA3_34
(
    .a(1'b1),
    .b(p11[32]),
    .s(CSA3_s[34]),
    .co(CSA3_co[34])
);

//CSA4
fa CSA4_0
(
    .a(p12[2]),
    .b(p13[0]),
    .c(y[27]),
    .s(CSA4_s[0]),
    .co(CSA4_co[0])
);
ha CSA4_1
(
    .a(p12[3]),
    .b(p13[1]),
    .s(CSA4_s[1]),
    .co(CSA4_co[1])
);
fa CSA4_2
(
    .a(p12[4]),
    .b(p13[2]),
    .c(p14[0]),
    .s(CSA4_s[2]),
    .co(CSA4_co[2])
);
fa CSA4_3
(
    .a(p12[5]),
    .b(p13[3]),
    .c(p14[1]),
    .s(CSA4_s[3]),
    .co(CSA4_co[3])
);
fa CSA4_4
(
    .a(p12[6]),
    .b(p13[4]),
    .c(p14[2]),
    .s(CSA4_s[4]),
    .co(CSA4_co[4])
);
fa CSA4_5
(
    .a(p12[7]),
    .b(p13[5]),
    .c(p14[3]),
    .s(CSA4_s[5]),
    .co(CSA4_co[5])
);
fa CSA4_6
(
    .a(p12[8]),
    .b(p13[6]),
    .c(p14[4]),
    .s(CSA4_s[6]),
    .co(CSA4_co[6])
);
fa CSA4_7
(
    .a(p12[9]),
    .b(p13[7]),
    .c(p14[5]),
    .s(CSA4_s[7]),
    .co(CSA4_co[7])
);
fa CSA4_8
(
    .a(p12[10]),
    .b(p13[8]),
    .c(p14[6]),
    .s(CSA4_s[8]),
    .co(CSA4_co[8])
);
fa CSA4_9
(
    .a(p12[11]),
    .b(p13[9]),
    .c(p14[7]),
    .s(CSA4_s[9]),
    .co(CSA4_co[9])
);
fa CSA4_10
(
    .a(p12[12]),
    .b(p13[10]),
    .c(p14[8]),
    .s(CSA4_s[10]),
    .co(CSA4_co[10])
);
fa CSA4_11
(
    .a(p12[13]),
    .b(p13[11]),
    .c(p14[9]),
    .s(CSA4_s[11]),
    .co(CSA4_co[11])
);
fa CSA4_12
(
    .a(p12[14]),
    .b(p13[12]),
    .c(p14[10]),
    .s(CSA4_s[12]),
    .co(CSA4_co[12])
);
fa CSA4_13
(
    .a(p12[15]),
    .b(p13[13]),
    .c(p14[11]),
    .s(CSA4_s[13]),
    .co(CSA4_co[13])
);
fa CSA4_14
(
    .a(p12[16]),
    .b(p13[14]),
    .c(p14[12]),
    .s(CSA4_s[14]),
    .co(CSA4_co[14])
);
fa CSA4_15
(
    .a(p12[17]),
    .b(p13[15]),
    .c(p14[13]),
    .s(CSA4_s[15]),
    .co(CSA4_co[15])
);
fa CSA4_16
(
    .a(p12[18]),
    .b(p13[16]),
    .c(p14[14]),
    .s(CSA4_s[16]),
    .co(CSA4_co[16])
);
fa CSA4_17
(
    .a(p12[19]),
    .b(p13[17]),
    .c(p14[15]),
    .s(CSA4_s[17]),
    .co(CSA4_co[17])
);
fa CSA4_18
(
    .a(p12[20]),
    .b(p13[18]),
    .c(p14[16]),
    .s(CSA4_s[18]),
    .co(CSA4_co[18])
);
fa CSA4_19
(
    .a(p12[21]),
    .b(p13[19]),
    .c(p14[17]),
    .s(CSA4_s[19]),
    .co(CSA4_co[19])
);
fa CSA4_20
(
    .a(p12[22]),
    .b(p13[20]),
    .c(p14[18]),
    .s(CSA4_s[20]),
    .co(CSA4_co[20])
);
fa CSA4_21
(
    .a(p12[23]),
    .b(p13[21]),
    .c(p14[19]),
    .s(CSA4_s[21]),
    .co(CSA4_co[21])
);
fa CSA4_22
(
    .a(p12[24]),
    .b(p13[22]),
    .c(p14[20]),
    .s(CSA4_s[22]),
    .co(CSA4_co[22])
);
fa CSA4_23
(
    .a(p12[25]),
    .b(p13[23]),
    .c(p14[21]),
    .s(CSA4_s[23]),
    .co(CSA4_co[23])
);
fa CSA4_24
(
    .a(p12[26]),
    .b(p13[24]),
    .c(p14[22]),
    .s(CSA4_s[24]),
    .co(CSA4_co[24])
);
fa CSA4_25
(
    .a(p12[27]),
    .b(p13[25]),
    .c(p14[23]),
    .s(CSA4_s[25]),
    .co(CSA4_co[25])
);
fa CSA4_26
(
    .a(p12[28]),
    .b(p13[26]),
    .c(p14[24]),
    .s(CSA4_s[26]),
    .co(CSA4_co[26])
);
fa CSA4_27
(
    .a(p12[29]),
    .b(p13[27]),
    .c(p14[25]),
    .s(CSA4_s[27]),
    .co(CSA4_co[27])
);
fa CSA4_28
(
    .a(p12[30]),
    .b(p13[28]),
    .c(p14[26]),
    .s(CSA4_s[28]),
    .co(CSA4_co[28])
);
fa CSA4_29
(
    .a(p12[31]),
    .b(p13[29]),
    .c(p14[27]),
    .s(CSA4_s[29]),
    .co(CSA4_co[29])
);
fa CSA4_30
(
    .a(p12[32]),
    .b(p13[30]),
    .c(p14[28]),
    .s(CSA4_s[30]),
    .co(CSA4_co[30])
);
fa CSA4_31
(
    .a(E[12]),
    .b(p13[31]),
    .c(p14[29]),
    .s(CSA4_s[31]),
    .co(CSA4_co[31])
);
fa CSA4_32
(
    .a(1'b1),
    .b(p13[32]),
    .c(p14[30]),
    .s(CSA4_s[32]),
    .co(CSA4_co[32])
);
ha CSA4_33
(
    .a(E[13]),
    .b(p14[31]),
    .s(CSA4_s[33]),
    .co(CSA4_co[33])
);
ha CSA4_34
(
    .a(1'b1),
    .b(p14[32]),
    .s(CSA4_s[34]),
    .co(CSA4_co[34])
);

//com
com_s com_0
(
    .a(CSA0_co[13]),
    .b(CSA1_co[7]),
    .c(CSA2_co[1]),
    .d(y[17]),
    .s(com_s[0]),
    .co(com_co[0]),
    .ca(com_ca[0])
);
fa com_1
(
    .a(CSA0_co[14]),
    .b(CSA1_co[8]),
    .c(CSA2_co[2]),
    .s(com_s[1]),
    .co(com_co[1])
);
com_s com_2
(
    .a(CSA0_co[15]),
    .b(CSA1_co[9]),
    .c(CSA2_co[3]),
    .d(p9[0]),
    .s(com_s[2]),
    .co(com_co[2]),
    .ca(com_ca[1])
);
com_s com_3
(
    .a(CSA0_co[16]),
    .b(CSA1_co[10]),
    .c(CSA2_co[4]),
    .d(p9[1]),
    .s(com_s[3]),
    .co(com_co[3]),
    .ca(com_ca[2])
);
fa com_4
(
    .a(CSA0_co[17]),
    .b(CSA1_co[11]),
    .c(CSA2_co[5]),
    .s(com_s[4]),
    .co(com_co[4])
);
com_s com_5
(
    .a(CSA0_co[18]),
    .b(CSA1_co[12]),
    .c(CSA2_co[6]),
    .d(CSA3_co[0]),
    .s(com_s[5]),
    .co(com_co[5]),
    .ca(com_ca[3])
);
com com_6
(
    .a(CSA0_co[19]),
    .b(CSA1_co[13]),
    .c(CSA2_co[7]),
    .d(CSA3_co[1]),
    .i(y[23]),
    .s(com_s[6]),
    .co(com_co[6]),
    .ca(com_ca[4])
);
com_s com_7
(
    .a(CSA0_co[20]),
    .b(CSA1_co[14]),
    .c(CSA2_co[8]),
    .d(CSA3_co[2]),
    .s(com_s[7]),
    .co(com_co[7]),
    .ca(com_ca[5])
);
com com_8
(
    .a(CSA0_co[21]),
    .b(CSA1_co[15]),
    .c(CSA2_co[9]),
    .d(CSA3_co[3]),
    .i(p12[0]),
    .s(com_s[8]),
    .co(com_co[8]),
    .ca(com_ca[6])
);
com com_9
(
    .a(CSA0_co[22]),
    .b(CSA1_co[16]),
    .c(CSA2_co[10]),
    .d(CSA3_co[4]),
    .i(p12[1]),
    .s(com_s[9]),
    .co(com_co[9]),
    .ca(com_ca[7])
);
com_s com_10
(
    .a(CSA0_co[23]),
    .b(CSA1_co[17]),
    .c(CSA2_co[11]),
    .d(CSA3_co[5]),
    .s(com_s[10]),
    .co(com_co[10]),
    .ca(com_ca[8])
);
com com_11
(
    .a(CSA0_co[24]),
    .b(CSA1_co[18]),
    .c(CSA2_co[12]),
    .d(CSA3_co[6]),
    .i(CSA4_co[0]),
    .s(com_s[11]),
    .co(com_co[11]),
    .ca(com_ca[9])
);
com com_12
(
    .a(CSA0_co[25]),
    .b(CSA1_co[19]),
    .c(CSA2_co[13]),
    .d(CSA3_co[7]),
    .i(CSA4_co[1]),
    .s(com_s[12]),
    .co(com_co[12]),
    .ca(com_ca[10])
);
com com_13
(
    .a(CSA0_co[26]),
    .b(CSA1_co[20]),
    .c(CSA2_co[14]),
    .d(CSA3_co[8]),
    .i(CSA4_co[2]),
    .s(com_s[13]),
    .co(com_co[13]),
    .ca(com_ca[11])
);
com com_14
(
    .a(CSA0_co[27]),
    .b(CSA1_co[21]),
    .c(CSA2_co[15]),
    .d(CSA3_co[9]),
    .i(CSA4_co[3]),
    .s(com_s[14]),
    .co(com_co[14]),
    .ca(com_ca[12])
);
com com_15
(
    .a(CSA0_co[28]),
    .b(CSA1_co[22]),
    .c(CSA2_co[16]),
    .d(CSA3_co[10]),
    .i(CSA4_co[4]),
    .s(com_s[15]),
    .co(com_co[15]),
    .ca(com_ca[13])
);
com com_16
(
    .a(CSA0_co[29]),
    .b(CSA1_co[23]),
    .c(CSA2_co[17]),
    .d(CSA3_co[11]),
    .i(CSA4_co[5]),
    .s(com_s[16]),
    .co(com_co[16]),
    .ca(com_ca[14])
);
com com_17
(
    .a(CSA0_co[30]),
    .b(CSA1_co[24]),
    .c(CSA2_co[18]),
    .d(CSA3_co[12]),
    .i(CSA4_co[6]),
    .s(com_s[17]),
    .co(com_co[17]),
    .ca(com_ca[15])
);
com com_18
(
    .a(CSA0_co[31]),
    .b(CSA1_co[25]),
    .c(CSA2_co[19]),
    .d(CSA3_co[13]),
    .i(CSA4_co[7]),
    .s(com_s[18]),
    .co(com_co[18]),
    .ca(com_ca[16])
);
com com_19
(
    .a(CSA0_co[32]),
    .b(CSA1_co[26]),
    .c(CSA2_co[20]),
    .d(CSA3_co[14]),
    .i(CSA4_co[8]),
    .s(com_s[19]),
    .co(com_co[19]),
    .ca(com_ca[17])
);
com com_20
(
    .a(CSA0_co[33]),
    .b(CSA1_co[27]),
    .c(CSA2_co[21]),
    .d(CSA3_co[15]),
    .i(CSA4_co[9]),
    .s(com_s[20]),
    .co(com_co[20]),
    .ca(com_ca[18])
);
com com_21
(
    .a(CSA0_co[34]),
    .b(CSA1_co[28]),
    .c(CSA2_co[22]),
    .d(CSA3_co[16]),
    .i(CSA4_co[10]),
    .s(com_s[21]),
    .co(com_co[21]),
    .ca(com_ca[19])
);
com_s com_22
(
    .a(CSA1_co[29]),
    .b(CSA2_co[23]),
    .c(CSA3_co[17]),
    .d(CSA4_co[11]),
    .s(com_s[22]),
    .co(com_co[22]),
    .ca(com_ca[20])
);
com_s com_23
(
    .a(CSA1_co[30]),
    .b(CSA2_co[24]),
    .c(CSA3_co[18]),
    .d(CSA4_co[12]),
    .s(com_s[23]),
    .co(com_co[23]),
    .ca(com_ca[21])
);
com_s com_24
(
    .a(CSA1_co[31]),
    .b(CSA2_co[25]),
    .c(CSA3_co[19]),
    .d(CSA4_co[13]),
    .s(com_s[24]),
    .co(com_co[24]),
    .ca(com_ca[22])
);
com_s com_25
(
    .a(CSA1_co[32]),
    .b(CSA2_co[26]),
    .c(CSA3_co[20]),
    .d(CSA4_co[14]),
    .s(com_s[25]),
    .co(com_co[25]),
    .ca(com_ca[23])
);
com_s com_26
(
    .a(CSA1_co[33]),
    .b(CSA2_co[27]),
    .c(CSA3_co[21]),
    .d(CSA4_co[15]),
    .s(com_s[26]),
    .co(com_co[26]),
    .ca(com_ca[24])
);
com_s com_27
(
    .a(CSA1_co[34]),
    .b(CSA2_co[28]),
    .c(CSA3_co[22]),
    .d(CSA4_co[16]),
    .s(com_s[27]),
    .co(com_co[27]),
    .ca(com_ca[25])
);
fa com_28
(
    .a(CSA2_co[29]),
    .b(CSA3_co[23]),
    .c(CSA4_co[17]),
    .s(com_s[28]),
    .co(com_co[28])
);
fa com_29
(
    .a(CSA2_co[30]),
    .b(CSA3_co[24]),
    .c(CSA4_co[18]),
    .s(com_s[29]),
    .co(com_co[29])
);
fa com_30
(
    .a(CSA2_co[31]),
    .b(CSA3_co[25]),
    .c(CSA4_co[19]),
    .s(com_s[30]),
    .co(com_co[30])
);
fa com_31
(
    .a(CSA2_co[32]),
    .b(CSA3_co[26]),
    .c(CSA4_co[20]),
    .s(com_s[31]),
    .co(com_co[31])
);
fa com_32
(
    .a(CSA2_co[33]),
    .b(CSA3_co[27]),
    .c(CSA4_co[21]),
    .s(com_s[32]),
    .co(com_co[32])
);
fa com_33
(
    .a(CSA2_co[34]),
    .b(CSA3_co[28]),
    .c(CSA4_co[21]),
    .s(com_s[33]),
    .co(com_co[33])
);


//CSA5
fa CSA5_0
(
    .a(CSA0_s[26]),
    .b(CSA1_s[20]),
    .c(y[29]),
    .s(CSA5_s[0]),
    .co(CSA5_co[0])
);
ha CSA5_1
(
    .a(CSA0_s[27]),
    .b(CSA1_s[21]),
    .s(CSA5_s[1]),
    .co(CSA5_co[1])
);
fa CSA5_2
(
    .a(CSA0_s[28]),
    .b(CSA1_s[22]),
    .c(p15[0]),
    .s(CSA5_s[2]),
    .co(CSA5_co[2])
);
fa CSA5_3
(
    .a(CSA0_s[29]),
    .b(CSA1_s[23]),
    .c(p15[1]),
    .s(CSA5_s[3]),
    .co(CSA5_co[3])
);
fa CSA5_4
(
    .a(CSA0_s[30]),
    .b(CSA1_s[24]),
    .c(p15[2]),
    .s(CSA5_s[4]),
    .co(CSA5_co[4])
);
fa CSA5_5
(
    .a(CSA0_s[31]),
    .b(CSA1_s[25]),
    .c(p15[3]),
    .s(CSA5_s[5]),
    .co(CSA5_co[5])
);
fa CSA5_6
(
    .a(CSA0_s[32]),
    .b(CSA1_s[26]),
    .c(p15[4]),
    .s(CSA5_s[6]),
    .co(CSA5_co[6])
);
fa CSA5_7
(
    .a(CSA0_s[33]),
    .b(CSA1_s[27]),
    .c(p15[5]),
    .s(CSA5_s[7]),
    .co(CSA5_co[7])
);
fa CSA5_8
(
    .a(CSA0_s[34]),
    .b(CSA1_s[28]),
    .c(p15[6]),
    .s(CSA5_s[8]),
    .co(CSA5_co[8])
);
fa CSA5_9
(
    .a(E[2]),
    .b(CSA1_s[29]),
    .c(p15[7]),
    .s(CSA5_s[9]),
    .co(CSA5_co[9])
);
fa CSA5_10
(
    .a(1'b1),
    .b(CSA1_s[30]),
    .c(p15[8]),
    .s(CSA5_s[10]),
    .co(CSA5_co[10])
);
ha CSA5_11
(
    .a(CSA1_s[31]),
    .b(p15[9]),
    .s(CSA5_s[11]),
    .co(CSA5_co[11])
);
ha CSA5_12
(
    .a(CSA1_s[32]),
    .b(p15[10]),
    .s(CSA5_s[12]),
    .co(CSA5_co[12])
);
ha CSA5_13
(
    .a(CSA1_s[33]),
    .b(p15[11]),
    .s(CSA5_s[13]),
    .co(CSA5_co[13])
);
ha CSA5_14
(
    .a(CSA1_s[34]),
    .b(p15[12]),
    .s(CSA5_s[14]),
    .co(CSA5_co[14])
);
ha CSA5_15
(
    .a(E[5]),
    .b(p15[13]),
    .s(CSA5_s[15]),
    .co(CSA5_co[15])
);
ha CSA5_16
(
    .a(1'b1),
    .b(p15[14]),
    .s(CSA5_s[16]),
    .co(CSA5_co[16])
);

//CSA6
fa CSA6_0
(
    .a(CSA2_s[10]),
    .b(CSA3_s[4]),
    .c(y[25]),
    .s(CSA6_s[0]),
    .co(CSA6_co[0])
);
ha CSA6_1
(
    .a(CSA2_s[11]),
    .b(CSA3_s[5]),
    .s(CSA6_s[1]),
    .co(CSA6_co[1])
);
generate
    genvar i;
    for(i = 2; i < 25 ;i = i + 1) 
    begin: g1
        fa CSA6_
        (
            .a(CSA2_s[i + 10]),
            .b(CSA3_s[i + 4]),
            .c(CSA4_s[i - 2]),
            .s(CSA6_s[i]),
            .co(CSA6_co[i])
        );
    end
endgenerate
fa CSA6_25
(
    .a(E[8]),
    .b(CSA3_s[29]),
    .c(CSA4_s[23]),
    .s(CSA6_s[25]),
    .co(CSA6_co[25])
);
fa CSA6_26
(
    .a(1'b1),
    .b(CSA3_s[30]),
    .c(CSA4_s[24]),
    .s(CSA6_s[26]),
    .co(CSA6_co[26])
);
ha CSA6_27
(
    .a(CSA3_s[31]),
    .b(CSA4_s[25]),
    .s(CSA6_s[27]),
    .co(CSA6_co[27])
);
ha CSA6_28
(
    .a(CSA3_s[32]),
    .b(CSA4_s[26]),
    .s(CSA6_s[28]),
    .co(CSA6_co[28])
);
ha CSA6_29
(
    .a(CSA3_s[33]),
    .b(CSA4_s[27]),
    .s(CSA6_s[29]),
    .co(CSA6_co[29])
);
ha CSA6_30
(
    .a(CSA3_s[34]),
    .b(CSA4_s[28]),
    .s(CSA6_s[30]),
    .co(CSA6_co[30])
);
ha CSA6_31
(
    .a(E[11]),
    .b(CSA4_s[29]),
    .s(CSA6_s[31]),
    .co(CSA6_co[31])
);
ha CSA6_32
(
    .a(1'b1),
    .b(CSA4_s[30]),
    .s(CSA6_s[32]),
    .co(CSA6_co[32])
);

//CSA7
fa CSA7_0
(
    .a(CSA1_co[1]),
    .b(y[11]),
    .c(CSA1_s[2]),
    .s(CSA7_s[0]),
    .co(CSA7_co[0])
);
ha CSA7_1
(
    .a(CSA1_co[2]),
    .b(CSA1_s[3]),
    .s(CSA7_s[1]),
    .co(CSA7_co[1])
);
fa CSA7_2
(
    .a(CSA1_co[3]),
    .b(p6[0]),
    .c(CSA1_s[4]),
    .s(CSA7_s[2]),
    .co(CSA7_co[2])
);
fa CSA7_3
(
    .a(CSA1_co[4]),
    .b(p6[1]),
    .c(CSA1_s[5]),
    .s(CSA7_s[3]),
    .co(CSA7_co[3])
);
ha CSA7_4
(
    .a(CSA1_co[5]),
    .b(CSA1_s[6]),
    .s(CSA7_s[4]),
    .co(CSA7_co[4])
);
fa CSA7_5
(
    .a(CSA1_co[6]),
    .b(CSA2_co[0]),
    .c(CSA1_s[7]),
    .s(CSA7_s[5]),
    .co(CSA7_co[5])
);
fa CSA7_6
(
    .a(com_co[0]),
    .b(com_ca[0]),
    .c(CSA1_s[9]),
    .s(CSA7_s[6]),
    .co(CSA7_co[6])
);
ha CSA7_7
(
    .a(com_co[1]),
    .b(CSA1_s[10]),
    .s(CSA7_s[7]),
    .co(CSA7_co[7])
);
fa CSA7_8
(
    .a(com_co[2]),
    .b(com_ca[1]),
    .c(CSA1_s[11]),
    .s(CSA7_s[8]),
    .co(CSA7_co[8])
);
fa CSA7_9
(
    .a(com_co[3]),
    .b(com_ca[2]),
    .c(CSA1_s[12]),
    .s(CSA7_s[9]),
    .co(CSA7_co[9])
);
ha CSA7_10
(
    .a(com_co[4]),
    .b(CSA1_s[13]),
    .s(CSA7_s[10]),
    .co(CSA7_co[10])
);
generate
    genvar ia;
    for(ia = 11; ia < 17 ;ia = ia + 1) 
    begin: g2
        fa CSA7_
        (
            .a(com_co[ia - 6]),
            .b(com_ca[ia - 8]),
            .c(CSA1_s[ia + 3]),
            .s(CSA7_s[ia]),
            .co(CSA7_co[ia])
        );
    end
endgenerate
ha CSA7_17
(
    .a(com_co[11]),
    .b(com_ca[9]),
    .s(CSA7_s[17]),
    .co(CSA7_co[17])
);
generate
    genvar ib;
    for(ib = 18; ib < 34 ;ib = ib + 1) 
    begin: g3
        fa CSA7_
        (
            .a(com_co[ib - 6]),
            .b(com_ca[ib - 8]),
            .c(CSA5_co[ib - 18]),
            .s(CSA7_s[ib]),
            .co(CSA7_co[ib])
        );
    end
endgenerate
ha CSA7_34
(
    .a(com_co[28]),
    .b(CSA5_co[16]),
    .s(CSA7_s[34]),
    .co(CSA7_co[34])
);

//CSA8
fa CSA8_0
(
    .a(CSA0_co[3]),
    .b(y[7]),
    .c(CSA0_s[4]),
    .s(CSA8_s[0]),
    .co(CSA8_co[0])
);
ha CSA8_1
(
    .a(CSA0_co[4]),
    .b(CSA0_s[5]),
    .s(CSA8_s[1]),
    .co(CSA8_co[1])
);
fa CSA8_2
(
    .a(CSA0_co[5]),
    .b(CSA1_s[0]),
    .c(CSA0_s[6]),
    .s(CSA8_s[2]),
    .co(CSA8_co[2])
);
fa CSA8_3
(
    .a(CSA0_co[6]),
    .b(CSA1_s[1]),
    .c(CSA0_s[7]),
    .s(CSA8_s[3]),
    .co(CSA8_co[3])
);
ha CSA8_4
(
    .a(CSA0_co[7]),
    .b(CSA0_s[8]),
    .s(CSA8_s[4]),
    .co(CSA8_co[4])
);
generate
    genvar ic;
    for(ic = 5; ic < 10 ;ic = ic + 1) 
    begin: g4
        fa CSA8_
        (
            .a(CSA0_co[ic + 3]),
            .b(CSA7_co[ic - 5]),
            .c(CSA0_s[ic + 4]),
            .s(CSA8_s[ic]),
            .co(CSA8_co[ic])
        );
    end
endgenerate
fa CSA8_10
(
    .a(com_s[0]),
    .b(CSA7_co[5]),
    .c(CSA0_s[14]),
    .s(CSA8_s[10]),
    .co(CSA8_co[10])
);
ha CSA8_11
(
    .a(com_s[1]),
    .b(CSA0_s[15]),
    .s(CSA8_s[11]),
    .co(CSA8_co[11])
);
generate
    genvar id;
    for(id = 12; id < 22 ;id = id + 1) 
    begin: g5
        fa CSA8_
        (
            .a(com_s[id - 10]),
            .b(CSA7_co[id - 6]),
            .c(CSA0_s[id + 4]),
            .s(CSA8_s[id]),
            .co(CSA8_co[id])
        );
    end
endgenerate
generate
    genvar ie;
    for(ie = 22; ie <  39;ie = ie + 1) 
    begin: g6
        fa CSA8_
        (
            .a(com_s[ie - 10]),
            .b(CSA7_co[ie - 6]),
            .c(CSA5_s[ie - 22]),
            .s(CSA8_s[ie]),
            .co(CSA8_co[ie])
        );
    end
endgenerate
fa CSA8_39
(
    .a(com_s[29]),
    .b(CSA7_co[33]),
    .c(p15[15]),
    .s(CSA8_s[39]),
    .co(CSA8_co[39])
);
fa CSA8_40
(
    .a(com_s[30]),
    .b(CSA7_co[34]),
    .c(p15[16]),
    .s(CSA8_s[40]),
    .co(CSA8_co[40])
);
generate
    genvar ig;
    for(ig = 41; ig <  44;ig = ig + 1) 
    begin: g7
        fa CSA8_
        (
            .a(com_s[ig - 10]),
            .b(com_co[ig - 11]),
            .c(p15[ig - 24]),
            .s(CSA8_s[ig]),
            .co(CSA8_co[ig])
        );
    end
endgenerate
fa CSA8_44
(
    .a(CSA3_co[29]),
    .b(com_co[33]),
    .c(p15[20]),
    .s(CSA8_s[44]),
    .co(CSA8_co[44])
);
generate
    genvar ih;
    for(ih = 45; ih <  50;ih = ih + 1) 
    begin: g8
        ha CSA8_
        (
            .a(CSA3_co[ih - 15]),
            .b(p15[ih - 24]),
            .s(CSA8_s[ih]),
            .co(CSA8_co[ih])
        );
    end
endgenerate

//CSA9
fa CSA9_0
(
    .a(CSA6_s[6]),
    .b(CSA6_co[5]),
    .c(y[31]),
    .s(CSA9_s[0]),
    .co(CSA9_co[0])
);
generate
    genvar ii;
    for(ii = 1; ii <  27; ii = ii + 1) 
    begin: g9
        ha CSA9_
        (
            .a(CSA6_s[ii + 6]),
            .b(CSA6_co[ii + 5]),
            .s(CSA9_s[ii]),
            .co(CSA9_co[ii])
        );
    end
endgenerate
ha CSA9_27
(
    .a(CSA4_s[31]),
    .b(CSA6_co[32]),
    .s(CSA9_s[27]),
    .co(CSA9_co[27])
);

//CSA10
fa CSA10_0
(
    .a(CSA8_co[5]),
    .b(CSA7_s[2]),
    .c(y[13]),
    .s(CSA10_s[0]),
    .co(CSA10_co[0])
);
ha CSA10_1
(
    .a(CSA8_co[6]),
    .b(CSA7_s[3]),
    .s(CSA10_s[1]),
    .co(CSA10_co[1])
);
fa CSA10_2
(
    .a(CSA8_co[7]),
    .b(CSA7_s[4]),
    .c(CSA2_s[0]),
    .s(CSA10_s[2]),
    .co(CSA10_co[2])
);
fa CSA10_3
(
    .a(CSA8_co[8]),
    .b(CSA7_s[5]),
    .c(CSA2_s[1]),
    .s(CSA10_s[3]),
    .co(CSA10_co[3])
);
fa CSA10_4
(
    .a(CSA8_co[9]),
    .b(CSA1_s[8]),
    .c(CSA2_s[2]),
    .s(CSA10_s[4]),
    .co(CSA10_co[4])
);
generate
    genvar ij;
    for(ij = 5; ij <  12; ij = ij + 1) 
    begin: g10
        fa CSA10_
        (
            .a(CSA8_co[ij + 5]),
            .b(CSA7_s[ij + 1]),
            .c(CSA2_s[ij - 2]),
            .s(CSA10_s[ij]),
            .co(CSA10_co[ij])
        );
    end
endgenerate
generate
    genvar ik;
    for(ik = 12; ik < 18; ik = ik + 1) 
    begin: g11
        fa CSA10_
        (
            .a(CSA8_co[ik + 5]),
            .b(CSA7_s[ik + 1]),
            .c(CSA6_s[ik - 12]),
            .s(CSA10_s[ik]),
            .co(CSA10_co[ik])
        );
    end
endgenerate
ha CSA10_18
(
    .a(CSA8_co[23]),
    .b(CSA7_s[19]),
    .s(CSA10_s[18]),
    .co(CSA10_co[18])
);
generate
    genvar il;
    for(il = 19; il < 34; il = il + 1) 
    begin: g12
        fa CSA10_
        (
            .a(CSA8_co[il + 5]),
            .b(CSA7_s[il + 1]),
            .c(CSA9_co[il - 19]),
            .s(CSA10_s[il]),
            .co(CSA10_co[il])
        );
    end
endgenerate
fa CSA10_34
(
    .a(CSA8_co[39]),
    .b(com_co[29]),
    .c(CSA9_co[15]),
    .s(CSA10_s[34]),
    .co(CSA10_co[34])
);
generate
    genvar im;
    for(im = 35; im < 38; im = im + 1) 
    begin: g13
        ha CSA10_
        (
            .a(CSA8_co[im + 5]),
            .b(CSA9_co[im - 19]),
            .s(CSA10_s[im]),
            .co(CSA10_co[im])
        );
    end
endgenerate
generate
    genvar in;
    for(in = 38; in < 45; in = in + 1) 
    begin: g14
        fa CSA10_
        (
            .a(CSA8_co[in + 5]),
            .b(CSA4_co[in - 15]),
            .c(CSA9_co[in - 19]),
            .s(CSA10_s[in]),
            .co(CSA10_co[in])
        );
    end
endgenerate
ha CSA10_45
(
    .a(CSA4_co[30]),
    .b(CSA9_co[26]),
    .s(CSA10_s[45]),
    .co(CSA10_co[45])
);
ha CSA10_46
(
    .a(CSA4_co[31]),
    .b(CSA9_co[27]),
    .s(CSA10_s[46]),
    .co(CSA10_co[46])
);


//CSA11
fa CSA11_0
(
    .a(CSA10_co[5]),
    .b(CSA8_s[12]),
    .c(y[19]),
    .s(CSA11_s[0]),
    .co(CSA11_co[0])
);
ha CSA11_1
(
    .a(CSA10_co[6]),
    .b(CSA8_s[13]),
    .s(CSA11_s[1]),
    .co(CSA11_co[1])
);
generate
    genvar io;
    for(io = 2; io < 6; io = io + 1) 
    begin: g15
        fa CSA11_
        (
            .a(CSA10_co[io + 5]),
            .b(CSA8_s[io + 12]),
            .c(CSA3_s[io - 2]),
            .s(CSA11_s[io]),
            .co(CSA11_co[io])
        );
    end
endgenerate
ha CSA11_6
(
    .a(CSA10_co[11]),
    .b(CSA8_s[18]),
    .s(CSA11_s[6]),
    .co(CSA11_co[6])
);
generate
    genvar ip;
    for(ip = 7; ip < 12; ip = ip + 1) 
    begin: g16
        fa CSA11_
        (
            .a(CSA10_co[ip + 5]),
            .b(CSA8_s[ip + 12]),
            .c(CSA6_co[ip - 7]),
            .s(CSA11_s[ip]),
            .co(CSA11_co[ip])
        );
    end
endgenerate
generate
    genvar iq;
    for(iq = 12; iq < 38; iq = iq + 1) 
    begin: g17
        fa CSA11_
        (
            .a(CSA10_co[iq + 5]),
            .b(CSA8_s[iq + 12]),
            .c(CSA9_s[iq - 12]),
            .s(CSA11_s[iq]),
            .co(CSA11_co[iq])
        );
    end
endgenerate
fa CSA11_38
(
    .a(CSA10_co[43]),
    .b(p15[26]),
    .c(CSA9_s[26]),
    .s(CSA11_s[38]),
    .co(CSA11_co[38])
);
fa CSA11_39
(
    .a(CSA10_co[44]),
    .b(p15[27]),
    .c(CSA9_s[27]),
    .s(CSA11_s[39]),
    .co(CSA11_co[39])
);
fa CSA11_40
(
    .a(CSA10_co[45]),
    .b(p15[28]),
    .c(CSA4_s[32]),
    .s(CSA11_s[40]),
    .co(CSA11_co[40])
);
fa CSA11_41
(
    .a(CSA10_co[46]),
    .b(p15[29]),
    .c(CSA4_s[33]),
    .s(CSA11_s[41]),
    .co(CSA11_co[41])
);
ha CSA11_42
(
    .a(p15[30]),
    .b(CSA4_s[34]),
    .s(CSA11_s[42]),
    .co(CSA11_co[42])
);
ha CSA11_43
(
    .a(p15[31]),
    .b(E[14]),
    .s(CSA11_s[43]),
    .co(CSA11_co[43])
);
ha CSA11_44
(
    .a(p15[32]),
    .b(1'b1),
    .s(CSA11_s[44]),
    .co(CSA11_co[44])
);

// CSA12
assign add0[0] = y[1];
assign add1[0] = p0[0];
assign add0[1] = 1'b0;
assign add1[1] = p0[1];
assign add0[2] = CSA0_s[0];
assign add1[2] = 1'b0;
assign add0[3] = CSA0_s[1];
assign add1[3] = CSA0_co[0];
assign add1[4] = 1'b0;

fa CSA12_4
(
    .a(CSA0_s[2]),
    .b(CSA0_co[1]),
    .c(y[5]),
    .s(add0[4]),
    .co(add1[5])
);
ha CSA12_5
(
    .a(CSA0_s[3]),
    .b(CSA0_co[2]),
    .s(add0[5]),
    .co(add1[6])
);
ha CSA12_6
(
    .a(CSA8_s[0]),
    .b(p3[0]),
    .s(add0[6]),
    .co(add1[7])
);
fa CSA12_7
(
    .a(CSA8_co[0]),
    .b(CSA8_s[1]),
    .c(p3[1]),
    .s(add0[7]),
    .co(add1[8])
);
ha CSA12_8
(
    .a(CSA8_co[1]),
    .b(CSA8_s[2]),
    .s(add0[8]),
    .co(add1[9])
);
fa CSA12_9
(
    .a(CSA8_co[2]),
    .b(CSA8_s[3]),
    .c(CSA1_co[0]),
    .s(add0[9]),
    .co(add1[10])
);
fa CSA12_10
(
    .a(CSA8_co[3]),
    .b(CSA8_s[4]),
    .c(CSA7_s[0]),
    .s(add0[10]),
    .co(add1[11])
);
fa CSA12_11
(
    .a(CSA8_co[4]),
    .b(CSA8_s[5]),
    .c(CSA7_s[1]),
    .s(add0[11]),
    .co(add1[12])
);
ha CSA12_12
(
    .a(CSA8_s[6]),
    .b(CSA10_s[0]),
    .s(add0[12]),
    .co(add1[13])
);
generate
    genvar ir;
    for(ir = 13; ir < 18; ir = ir + 1) 
    begin: g18
        fa CSA12_
        (
            .a(CSA10_co[ir - 13]),
            .b(CSA8_s[ir - 6]),
            .c(CSA10_s[ir - 12]),
            .s(add0[ir]),
            .co(add1[ir + 1])
        );
    end
endgenerate
ha CSA12_18
(
    .a(CSA11_s[0]),
    .b(CSA10_s[6]),
    .s(add0[18]),
    .co(add1[19])
);
generate
    genvar is;
    for(is = 19; is < 59; is = is + 1) 
    begin: g19
        fa CSA12_
        (
            .a(CSA11_co[is - 19]),
            .b(CSA11_s[is - 18]),
            .c(CSA10_s[is - 12]),
            .s(add0[is]),
            .co(add1[is + 1])
        );
    end
endgenerate
generate
    genvar it;
    for(it = 59; it < 62; it = it + 1) 
    begin: g20
        fa CSA12_
        (
            .a(CSA11_co[it - 19]),
            .b(CSA11_s[it - 18]),
            .c(CSA4_co[it - 27]),
            .s(add0[it]),
            .co(add1[it + 1])
        );
    end
endgenerate
ha CSA12_62
(
    .a(CSA11_co[43]),
    .b(CSA11_s[44]),
    .s(add0[62]),
    .co(add1[63])
);

assign add0[63] = CSA11_co[44] + E[15];


// //=======================================================
// wire [63:0] test11c;
// wire [63:0] test11s;
// wire [63:0] test10s;

// assign test11c[0] = y[1];
// assign test11c[1] = 0;
// assign test11c[5 : 2] = CSA0_s[3 : 0];
// assign test11c[6] = 0;
// assign test11c[11 : 7] = CSA8_co[4 : 0];
// assign test11c[12] = 0;
// assign test11c[17 : 13] = CSA10_co[4 : 0];
// assign test11c[18] = 0;
// assign test11c[63 : 19] = CSA11_co[44 : 0];

// assign test11s[1 : 0] = p0[1 : 0];
// assign test11s[2] = 0;
// assign test11s[5 : 3] = CSA0_co[2 : 0];
// assign test11s[17 : 6] = CSA8_s[11 : 0];
// assign test11s[62 : 18] = CSA11_s[44 : 0];
// assign test11s[63] = E[15];

// assign test10s[3 : 0] = 0;
// assign test10s[4] = y[5];
// assign test10s[5] = 0;
// assign test10s[7 : 6] = p3[1 : 0];
// assign test10s[8] = 0;
// assign test10s[9] = CSA1_co[0];
// assign test10s[11 : 10] = CSA7_s[1 : 0];
// assign test10s[58 : 12] = CSA10_s[46 : 0];
// assign test10s[61 : 59] = CSA4_co[34 : 32];
// assign test10s[63 : 62] = 0;

// wire [63 : 0] test0s;
// wire [63 : 0] test0c;
// wire [63 : 0] test1s;
// wire [63 : 0] test1c;
// wire [63 : 0] test2s;
// wire [63 : 0] test2c;
// wire [63 : 0] test3s;
// wire [63 : 0] test3c;
// wire [63 : 0] test4s;
// wire [63 : 0] test4c;

// wire [63 : 0] test0;
// wire [63 : 0] test1;
// wire [63 : 0] test2;
// wire [63 : 0] test3;
// wire [63 : 0] test4;
// wire [63 : 0] test5;
// wire [63 : 0] test6;
// wire [63 : 0] test7;
// wire [63 : 0] test8;
// wire [63 : 0] test9;
// wire [63 : 0] test10;
// wire [63 : 0] test11;
// wire [63 : 0] test12;
// wire [63 : 0] test13;
// wire [63 : 0] test14;
// wire [63 : 0] test15;
// wire [63 : 0] test16;

// assign test0c[1 : 0] = p0[1 : 0];
// assign test0c[2] = 0;
// assign test0c[37 : 3] = CSA0_co[34 : 0];
// assign test0c[63 : 38] = 0;

// assign test0s[0] = y[1];
// assign test0s[1] = 0;
// assign test0s[36 : 2] = CSA0_s[34 : 0];
// assign test0s[37] = E[2];
// assign test0s[38] = 1;
// assign test0s[63 : 39] = 0;

// assign test1c[3 : 0] = 0;
// assign test1c[4] = y[5];
// assign test1c[5] = 0;
// assign test1c[7 : 6] = p3[1 : 0];
// assign test1c[8] = 0;
// assign test1c[43 : 9] = CSA1_co[34 : 0];
// assign test1c[63 : 44] = 0;

// assign test1s[5 : 0] = 0;
// assign test1s[6] = y[7];
// assign test1s[7] = 0;
// assign test1s[42 : 8] = CSA1_s[34 : 0];
// assign test1s[43] = E[5];
// assign test1s[44] = 1;
// assign test1s[63 : 45] = 0;

// assign test2c[9 : 0] = 0;
// assign test2c[10] = y[11];
// assign test2c[11] = 0;
// assign test2c[13 : 12] = p6[1 : 0];
// assign test2c[14] = 0;
// assign test2c[49 : 15] = CSA2_co[34 : 0];
// assign test2c[63 : 50] = 0;

// assign test2s[11 : 0] = 0;
// assign test2s[12] = y[13];
// assign test2s[13] = 0;
// assign test2s[48 : 14] = CSA2_s[34 : 0];
// assign test2s[49] = E[8];
// assign test2s[50] = 1;
// assign test2s[63 : 51] = 0;


// assign test3c[15 : 0] = 0;
// assign test3c[16] = y[17];
// assign test3c[17] = 0;
// assign test3c[19 : 18] = p9[1 : 0];
// assign test3c[20] = 0;
// assign test3c[55 : 21] = CSA3_co[34 : 0];
// assign test3c[63 : 56] = 0;

// assign test3s[17 : 0] = 0;
// assign test3s[18] = y[19];
// assign test3s[19] = 0;
// assign test3s[54 : 20] = CSA3_s[34 : 0];
// assign test3s[55] = E[11];
// assign test3s[56] = 1;
// assign test3s[63 : 57] = 0;

// assign test4c[21 : 0] = 0;
// assign test4c[22] = y[23];
// assign test4c[23] = 0;
// assign test4c[25 : 24] = p12[1 : 0];
// assign test4c[26] = 0;
// assign test4c[61 : 27] = CSA4_co[34 : 0];
// assign test4c[63 : 62] = 0;

// assign test4s[23 : 0] = 0;
// assign test4s[24] = y[25];
// assign test4s[25] = 0;
// assign test4s[60 : 26] = CSA4_s[34 : 0];
// assign test4s[61] = E[14];
// assign test4s[62] = 1;
// assign test4s[63] = 0;

// assign test0[32 : 0] = p0[32 : 0];
// assign test0[33] = ~E[0];
// assign test0[34] = ~E[0];
// assign test0[63 : 35] = E[0];

// assign test1[0] = y[1];
// assign test1[1] = 0;
// assign test1[34 : 2] = p1[32 : 0];
// assign test1[35] = E[1];
// assign test1[36] = 1;
// assign test1[63 : 37] = 0;

// assign test2[1 : 0] = 0;
// assign test2[2] = y[3];
// assign test2[3] = 0;
// assign test2[36 : 4] = p2[32 : 0];
// assign test2[37] = E[2];
// assign test2[38] = 1;
// assign test2[63 : 39] = 0;

// assign test3[3 : 0] = 0;
// assign test3[4] = y[5];
// assign test3[5] = 0;
// assign test3[38 : 6] = p3[32 : 0];
// assign test3[39] = E[3];
// assign test3[40] = 1;
// assign test3[63 : 41] = 0;


// assign test4[5 : 0] = 0;
// assign test4[6] = y[7];
// assign test4[7] = 0;
// assign test4[40 : 8] = p4[32 : 0];
// assign test4[41] = E[4];
// assign test4[42] = 1;
// assign test4[63 : 43] = 0;

// assign test5[7 : 0] = 0;
// assign test5[8] = y[9];
// assign test5[9] = 0;
// assign test5[42 : 10] = p5[32 : 0];
// assign test5[43] = E[5];
// assign test5[44] = 1;
// assign test5[63 : 45] = 0;

// assign test6[9 : 0] = 0;
// assign test6[10] = y[11];
// assign test6[11] = 0;
// assign test6[44 : 12] = p6[32 : 0];
// assign test6[45] = E[6];
// assign test6[46] = 1;
// assign test6[63 : 47] = 0;

// assign test7[11 : 0] = 0;
// assign test7[12] = y[13];
// assign test7[13] = 0;
// assign test7[46 : 14] = p7[32 : 0];
// assign test7[47] = E[7];
// assign test7[48] = 1;
// assign test7[63 : 49] = 0;

// assign test8[13 : 0] = 0;
// assign test8[14] = y[15];
// assign test8[15] = 0;
// assign test8[48 : 16] = p8[32 : 0];
// assign test8[49] = E[8];
// assign test8[50] = 1;
// assign test8[63 : 51] = 0;

// assign test9[15 : 0] = 0;
// assign test9[16] = y[17];
// assign test9[17] = 0;
// assign test9[50 : 18] = p9[32 : 0];
// assign test9[51] = E[9];
// assign test9[52] = 1;
// assign test9[63 : 53] = 0;

// assign test10[17 : 0] = 0;
// assign test10[18] = y[19];
// assign test10[19] = 0;
// assign test10[52 : 20] = p10[32 : 0];
// assign test10[53] = E[10];
// assign test10[54] = 1;
// assign test10[63 : 55] = 0;

// assign test11[19 : 0] = 0;
// assign test11[20] = y[21];
// assign test11[21] = 0;
// assign test11[54 : 22] = p11[32 : 0];
// assign test11[55] = E[11];
// assign test11[56] = 1;
// assign test11[63 : 57] = 0;

// assign test12[21 : 0] = 0;
// assign test12[22] = y[23];
// assign test12[23] = 0;
// assign test12[56 : 24] = p12[32 : 0];
// assign test12[57] = E[12];
// assign test12[58] = 1;
// assign test12[63 : 59] = 0;

// assign test13[23 : 0] = 0;
// assign test13[24] = y[25];
// assign test13[25] = 0;
// assign test13[58 : 26] = p13[32 : 0];
// assign test13[59] = E[13];
// assign test13[60] = 1;
// assign test13[63 : 61] = 0;

// assign test14[25 : 0] = 0;
// assign test14[26] = y[27];
// assign test14[27] = 0;
// assign test14[60 : 28] = p13[32 : 0];
// assign test14[61] = E[14];
// assign test14[62] = 1;
// assign test14[63] = 0;


// assign test15[27 : 0] = 0;
// assign test15[28] = y[29];
// assign test15[29] = 0;
// assign test15[62 : 30] = p15[32 : 0];
// assign test15[63] = E[15];

// assign test16[29 : 0] = 0;
// assign test16[30] = y[31];
// assign test16[63 : 31] = 0;

// assign add0 = test4c + test4s;
// assign add1 = test3c + test3s + test2c + test2s + test1c + test1s + test0c + test0s + test15 + test16;

// // assign add0 = 0;
// // assign add1 = test0 + test1 + test2 +test3 +test4 +test5 +test6 +test7 +test8 +test9 +test10 +test11 +test12 +test13 +test14 +test15 +test16;


endmodule